-- probe.vhd

-- Generated using ACDS version 21.1 850

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity probe is
	port (
		probe : in std_logic_vector(95 downto 0) := (others => '0')  -- probes.probe
	);
end entity probe;

architecture rtl of probe is
	component altsource_probe_top is
		generic (
			sld_auto_instance_index : string  := "YES";
			sld_instance_index      : integer := 0;
			instance_id             : string  := "NONE";
			probe_width             : integer := 1;
			source_width            : integer := 1;
			enable_metastability    : string  := "NO"
		);
		port (
			probe : in std_logic_vector(95 downto 0) := (others => 'X')  -- probe
		);
	end component altsource_probe_top;

begin

	in_system_sources_probes_0 : component altsource_probe_top
		generic map (
			sld_auto_instance_index => "YES",
			sld_instance_index      => 0,
			instance_id             => "NONE",
			probe_width             => 96,
			source_width            => 0,
			enable_metastability    => "NO"
		)
		port map (
			probe => probe  -- probes.probe
		);

end architecture rtl; -- of probe
