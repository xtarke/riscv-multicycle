-------------------------------------------------------------------
-- Name        : de0_lite.vhd
-- Author      : 
-- Version     : 0.1
-- Copyright   : Departamento de Eletrônica, Florianópolis, IFSC
-- Description : Projeto base DE10-Lite
-------------------------------------------------------------------
LIBRARY ieee;
USE IEEE.STD_LOGIC_1164.ALL;

entity de0_lite is 
	port (
		---------- CLOCK ----------
		ADC_CLK_10:	in std_logic;
		MAX10_CLK1_50: in std_logic;
		MAX10_CLK2_50: in std_logic;
		
		----------- SDRAM ------------
		DRAM_ADDR: out std_logic_vector (12 downto 0);
		DRAM_BA: out std_logic_vector (1 downto 0);
		DRAM_CAS_N: out std_logic;
		DRAM_CKE: out std_logic;
		DRAM_CLK: out std_logic;
		DRAM_CS_N: out std_logic;		
		DRAM_DQ: inout std_logic_vector(15 downto 0);
		DRAM_LDQM: out std_logic;
		DRAM_RAS_N: out std_logic;
		DRAM_UDQM: out std_logic;
		DRAM_WE_N: out std_logic;
		
		----------- SEG7 ------------
		HEX0: out std_logic_vector(7 downto 0);
		HEX1: out std_logic_vector(7 downto 0);
		HEX2: out std_logic_vector(7 downto 0);
		HEX3: out std_logic_vector(7 downto 0);
		HEX4: out std_logic_vector(7 downto 0);
		HEX5: out std_logic_vector(7 downto 0);

		----------- KEY ------------
		KEY: in std_logic_vector(1 downto 0);

		----------- LED ------------
		LEDR: out std_logic_vector(9 downto 0);

		----------- SW ------------
		SW: in std_logic_vector(9 downto 0);

		----------- VGA ------------
		VGA_B: out std_logic_vector(3 downto 0);
		VGA_G: out std_logic_vector(3 downto 0);
		VGA_HS: out std_logic;
		VGA_R: out std_logic_vector(3 downto 0);
		VGA_VS: out std_logic;
	
		----------- Accelerometer ------------
		GSENSOR_CS_N: out std_logic;
		GSENSOR_INT: in std_logic_vector(2 downto 1);
		GSENSOR_SCLK: out std_logic;
		GSENSOR_SDI: inout std_logic;
		GSENSOR_SDO: inout std_logic;
	
		----------- Arduino ------------
		ARDUINO_IO: inout std_logic_vector(15 downto 0);
		ARDUINO_RESET_N: inout std_logic
	);
end entity;


architecture rtl of de0_lite is
	signal clock : std_logic;
	signal clock2 : std_logic  := '0';
	signal jmp   : std_logic;
	signal counter : integer  :=  0;
	signal inp : std_logic;
	signal div : integer range 0 to 50;
	
begin
	
	pll: ENTITY work.pll_500khz 
	PORT map
	(
		inclk0	 => MAX10_CLK1_50,
		c0		 => clock
	);
	
	spi: entity work.SPI
	port map(
	  i_clk  	 => clock,                   
	  i_rst      => SW(9),        
	  i_tx_start => KEY(1),         
	  i_data     => SW(7 downto 0),        
	  i_miso     => ARDUINO_IO(4),        
	  o_data     => LEDR(7 downto 0),      
	  o_tx_end   => ARDUINO_IO(0),       
	  o_sclk     => ARDUINO_IO(1),       
	  o_ss       => ARDUINO_IO(2),      
	  o_mosi     => ARDUINO_IO(3),
	  debug_idle_flag  => ARDUINO_IO(5),
	  debug_tx_flag    => ARDUINO_IO(6),
	  debug_end_flag   => ARDUINO_IO(7)      
	);
	
--	process(clock)
--	begin
--		if rising_edge(clock) then
--			div  <=  div +1;
--			if div = 0 then
--				clock2  <=  not clock2;
--			end if;
--		end if;
--	end process;
	
--	process(clock,KEY(1))
--	begin
--		if rising_edge(clock) and KEY(1) = '1' then
--			counter  <=  counter + 1;
--			inp  <= '1';
--			
--			if counter <= 32 then
--				inp  <= '0';
--			end if;
--		end if;
--		if KEY(1) = '0' then	
--			counter  <= 0;
--		end if;
--		
--	end process;
end;

