// TODO "Go back"
//      Navigate back to `step_2_navigation` by pressing **Alt+Left key**
`ifndef _constants_svh_
`define _constants_svh_

`define MAX_COUNT 2 ** 8 - 1

`define ANSWER 4 * 10 + 2

`define MAGIC_NUMBER 16'hda01

`endif
