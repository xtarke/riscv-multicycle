
module probe (
	probe);	

	input	[95:0]	probe;
endmodule
