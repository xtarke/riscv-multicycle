-------------------------------------------------------------------
-- Name        : de0_lite.vhd
-- Author      : 
-- Version     : 0.1
-- Copyright   : Departamento de Eletrônica, Florianópolis, IFSC
-- Description : Projeto base DE10-Lite
-------------------------------------------------------------------
LIBRARY ieee;
USE IEEE.STD_LOGIC_1164.ALL;

entity de10_lite is 
	port (
		---------- CLOCK ----------
		ADC_CLK_10:	in std_logic;
		MAX10_CLK1_50: in std_logic;
		MAX10_CLK2_50: in std_logic;
		
		----------- SDRAM ------------
		DRAM_ADDR: out std_logic_vector (12 downto 0);
		DRAM_BA: out std_logic_vector (1 downto 0);
		DRAM_CAS_N: out std_logic;
		DRAM_CKE: out std_logic;
		DRAM_CLK: out std_logic;
		DRAM_CS_N: out std_logic;		
		DRAM_DQ: inout std_logic_vector(15 downto 0);
		DRAM_LDQM: out std_logic;
		DRAM_RAS_N: out std_logic;
		DRAM_UDQM: out std_logic;
		DRAM_WE_N: out std_logic;
		
		----------- SEG7 ------------
		HEX0: out std_logic_vector(7 downto 0);
		HEX1: out std_logic_vector(7 downto 0);
		HEX2: out std_logic_vector(7 downto 0);
		HEX3: out std_logic_vector(7 downto 0);
		HEX4: out std_logic_vector(7 downto 0);
		HEX5: out std_logic_vector(7 downto 0);

		----------- KEY ------------
		KEY: in std_logic_vector(1 downto 0);

		----------- LED ------------
		LEDR: out std_logic_vector(9 downto 0);

		----------- SW ------------
		SW: in std_logic_vector(9 downto 0);

		----------- VGA ------------
		VGA_B: out std_logic_vector(3 downto 0);
		VGA_G: out std_logic_vector(3 downto 0);
		VGA_HS: out std_logic;
		VGA_R: out std_logic_vector(3 downto 0);
		VGA_VS: out std_logic;
	
		----------- Accelerometer ------------
		GSENSOR_CS_N: out std_logic;
		GSENSOR_INT: in std_logic_vector(2 downto 1);
		GSENSOR_SCLK: out std_logic;
		GSENSOR_SDI: inout std_logic;
		GSENSOR_SDO: inout std_logic;
	
		----------- Arduino ------------
		ARDUINO_IO: inout std_logic_vector(15 downto 0);
		ARDUINO_RESET_N: inout std_logic
	);
end entity;


architecture rtl of de10_lite is

		--source envia dados (write_data)
		--probe le dados (read_data)
		--component probes is
		--	port (
		--		source : out std_logic_vector(31 downto 0);                    -- source
		--		probe  : in  std_logic_vector(31 downto 0) := (others => 'X')  -- probe
		--	);
		--end component probes;
		
		--sinais do probes
		--signal probe : std_logic_vector(31 downto 0);
		--signal source : std_logic_vector(31 downto 0);
		
		--sinais do rng
		signal clk : std_logic;  -- clock do sistema
		signal rst : std_logic;  -- reset sincrono
      signal chip_select : std_logic; -- ativa este periferico
		signal addr : std_logic_vector(1 downto 0);  -- seleciona registrador
		signal read_data : std_logic_vector(31 downto 0); -- valor lido pelo CPU

	
begin

		--instacia IP probes
		--u0 : component probes
		--	port map (
		--		source => source,
		--		probe  => probe
		--	);

		--instancia IP rng
		dut_rng: entity work.rng
		  port map(
				clk         => SW(8),
				rst         => SW(9),
				chip_select  => SW(1),
				addr         => SW(3 downto 2),
				read_data    => read_data
		  );

		--instancia IP display
		dut0 : entity work.seven_seg
			port map (
				input  => read_data(3 downto 0), 
				output => HEX0
			);
			
		dut1 : entity work.seven_seg
			port map (
				input  => read_data(7 downto 4), 
				output => HEX1
			);
			
		dut2 : entity work.seven_seg
			port map (
				input  => read_data(11 downto 8), 
				output => HEX2
			);
			
		dut3 : entity work.seven_seg
			port map (
				input  => read_data(15 downto 12), 
				output => HEX3
			);
			
		dut4 : entity work.seven_seg
			port map (
				input  => read_data(19 downto 16), 
				output => HEX4
			);

		dut5 : entity work.seven_seg
			port map (
				input  => read_data(23 downto 20), 
				output => HEX5
			);
			
		--write_data <= std_logic_vector(source(31 downto 0)); --escrever nova seed
		--probe(31 downto 0) <= std_logic_vector(read_data(31 downto 0)); -- ler número gerado

end architecture;
