PLL_100KHz_inst : PLL_100KHz PORT MAP (
		inclk0	 => inclk0_sig,
		c0	 => c0_sig
	);
