library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity sram is
	port(
		clk : in std_logic;
		rst : in std_logic
	);
end entity sram;

architecture RTL of sram is
	
begin

end architecture RTL;
