library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity lookup_angle is
    port(
        raw_in    : in  std_logic_vector(7 downto 0); -- Entrada "crua" (0..255)
        signal_bit : in  STD_LOGIC; -- Sinal da entrada (0 = positivo, 1 = negativo)
        angle_out : out std_logic_vector(7 downto 0)  -- Ângulo correspondente (0..90)
    );
end entity lookup_angle;

architecture rtl of lookup_angle is
    -- Define um tipo de array para a LUT com entradas de 8 bits
    type lut_array is array (0 to 280) of std_logic_vector(7 downto 0);
    type neg_lut_array is array (0 to 270) of std_logic_vector(7 downto 0);

    -- Exemplo de tabela – preencha todos os valores conforme sua relação.
    constant angle_table : lut_array := (
        280 => "01011010",
        279 => "01011010",
        278 => "01011010",
        277 => "01011010",
        276 => "01011010",
        275 => "01011010",
        274 => "01011010",
        273 => "01011010",
        272 => "01011010",
        271 => "01011010",
        270 => "01011010",
        269 => "01011010",
        268 => "01011010",
        267 => "01011010",
        266 => "01011010",
        265 => "01011010",
        264 => "01011010",
        263 => "01011010",
        262 => "01011010",
        261 => "01011010",
        260 => "01011010",
        259 => "01011010",
        258 => "01011010",
        257 => "01011010",
        256 => "01011010",
        255 => "01011010",
        254 => "01010101",
        253 => "01010011",
        252 => "01010001",
        251 => "01010000",
        250 => "01001111",
        249 => "01001110",
        248 => "01001101",
        247 => "01001100",
        246 => "01001011",
        245 => "01001010",
        244 => "01001001",
        243 => "01001000",
        242 => "01001000",
        241 => "01000111",
        240 => "01000110",
        239 => "01000110",
        238 => "01000101",
        237 => "01000100",
        236 => "01000100",
        235 => "01000011",
        234 => "01000011",
        233 => "01000010",
        232 => "01000001",
        231 => "01000001",
        230 => "01000000",
        229 => "01000000",
        228 => "00111111",
        227 => "00111111",
        226 => "00111110",
        225 => "00111110",
        224 => "00111101",
        223 => "00111101",
        222 => "00111101",
        221 => "00111100",
        220 => "00111100",
        219 => "00111011",
        218 => "00111011",
        217 => "00111010",
        216 => "00111010",
        215 => "00111001",
        214 => "00111001",
        213 => "00111001",
        212 => "00111000",
        211 => "00111000",
        210 => "00110111",
        209 => "00110111",
        208 => "00110111",
        207 => "00110110",
        206 => "00110110",
        205 => "00110110",
        204 => "00110101",
        203 => "00110101",
        202 => "00110100",
        201 => "00110100",
        200 => "00110100",
        199 => "00110011",
        198 => "00110011",
        197 => "00110011",
        196 => "00110010",
        195 => "00110010",
        194 => "00110010",
        193 => "00110001",
        192 => "00110001",
        191 => "00110001",
        190 => "00110000",
        189 => "00110000",
        188 => "00101111",
        187 => "00101111",
        186 => "00101111",
        185 => "00101111",
        184 => "00101110",
        183 => "00101110",
        182 => "00101110",
        181 => "00101101",
        180 => "00101101",
        179 => "00101101",
        178 => "00101100",
        177 => "00101100",
        176 => "00101100",
        175 => "00101011",
        174 => "00101011",
        173 => "00101011",
        172 => "00101010",
        171 => "00101010",
        170 => "00101010",
        169 => "00101010",
        168 => "00101001",
        167 => "00101001",
        166 => "00101001",
        165 => "00101000",
        164 => "00101000",
        163 => "00101000",
        162 => "00100111",
        161 => "00100111",
        160 => "00100111",
        159 => "00100111",
        158 => "00100110",
        157 => "00100110",
        156 => "00100110",
        155 => "00100101",
        154 => "00100101",
        153 => "00100101",
        152 => "00100101",
        151 => "00100100",
        150 => "00100100",
        149 => "00100100",
        148 => "00100011",
        147 => "00100011",
        146 => "00100011",
        145 => "00100011",
        144 => "00100010",
        143 => "00100010",
        142 => "00100010",
        141 => "00100010",
        140 => "00100001",
        139 => "00100001",
        138 => "00100001",
        137 => "00100000",
        136 => "00100000",
        135 => "00100000",
        134 => "00100000",
        133 => "00011111",
        132 => "00011111",
        131 => "00011111",
        130 => "00011111",
        129 => "00011110",
        128 => "00011110",
        127 => "00011110",
        126 => "00011110",
        125 => "00011101",
        124 => "00011101",
        123 => "00011101",
        122 => "00011101",
        121 => "00011100",
        120 => "00011100",
        119 => "00011100",
        118 => "00011100",
        117 => "00011011",
        116 => "00011011",
        115 => "00011011",
        114 => "00011011",
        113 => "00011010",
        112 => "00011010",
        111 => "00011010",
        110 => "00011010",
        109 => "00011001",
        108 => "00011001",
        107 => "00011001",
        106 => "00011001",
        105 => "00011000",
        104 => "00011000",
        103 => "00011000",
        102 => "00011000",
        101 => "00010111",
        100 => "00010111",
        99 => "00010111",
        98 => "00010111",
        97 => "00010110",
        96 => "00010110",
        95 => "00010110",
        94 => "00010110",
        93 => "00010101",
        92 => "00010101",
        91 => "00010101",
        90 => "00010101",
        89 => "00010100",
        88 => "00010100",
        87 => "00010100",
        86 => "00010100",
        85 => "00010011",
        84 => "00010011",
        83 => "00010011",
        82 => "00010011",
        81 => "00010011",
        80 => "00010010",
        79 => "00010010",
        78 => "00010010",
        77 => "00010010",
        76 => "00010001",
        75 => "00010001",
        74 => "00010001",
        73 => "00010001",
        72 => "00010000",
        71 => "00010000",
        70 => "00010000",
        69 => "00010000",
        68 => "00001111",
        67 => "00001111",
        66 => "00001111",
        65 => "00001111",
        64 => "00001111",
        63 => "00001110",
        62 => "00001110",
        61 => "00001110",
        60 => "00001110",
        59 => "00001101",
        58 => "00001101",
        57 => "00001101",
        56 => "00001101",
        55 => "00001100",
        54 => "00001100",
        53 => "00001100",
        52 => "00001100",
        51 => "00001100",
        50 => "00001011",
        49 => "00001011",
        48 => "00001011",
        47 => "00001011",
        46 => "00001010",
        45 => "00001010",
        44 => "00001010",
        43 => "00001010",
        42 => "00001001",
        41 => "00001001",
        40 => "00001001",
        39 => "00001001",
        38 => "00001001",
        37 => "00001000",
        36 => "00001000",
        35 => "00001000",
        34 => "00001000",
        33 => "00000111",
        32 => "00000111",
        31 => "00000111",
        30 => "00000111",
        29 => "00000111",
        28 => "00000110",
        27 => "00000110",
        26 => "00000110",
        25 => "00000110",
        24 => "00000101",
        23 => "00000101",
        22 => "00000101",
        21 => "00000101",
        20 => "00000100",
        19 => "00000100",
        18 => "00000100",
        17 => "00000100",
        16 => "00000100",
        15 => "00000011",
        14 => "00000011",
        13 => "00000011",
        12 => "00000011",
        11 => "00000010",
        10 => "00000010",
        9 => "00000010",
        8 => "00000010",
        7 => "00000010",
        6 => "00000001",
        5 => "00000001",
        4 => "00000001",
        3 => "00000001",
        2 => "00000000",
        1 => "00000000",
        0 => "00000000"
    );
    
    constant negative_angle_table : neg_lut_array := (
        270 => "01011010",
        269 => "01011010",
        268 => "01011010",
        267 => "01011010",
        266 => "01011010",
        265 => "01011010",
        264 => "01011010",
        263 => "01011010",
        262 => "01011010",
        261 => "01011010",
        260 => "01011010",
        259 => "01011010",
        258 => "01011010",
        257 => "01011010",
        256 => "01011010",
        255 => "01011010",
        254 => "01011010",
        253 => "01011010",
        252 => "01011010",
        251 => "01011010",
        250 => "01011010",
        249 => "01011010",
        248 => "01011010",
        247 => "01011010",
        246 => "01011010",
        245 => "01011010",
        244 => "01011010",
        243 => "01011010",
        242 => "01011010",
        241 => "01011010",
        240 => "01011010",
        239 => "01011010",
        238 => "01011010",
        237 => "01011010",
        236 => "01011010",
        235 => "01011010",
        234 => "01011010",
        233 => "01011010",
        232 => "01011010",
        231 => "01011010",
        230 => "01011010",
        229 => "01010101",
        228 => "01010010",
        227 => "01010001",
        226 => "01001111",
        225 => "01001110",
        224 => "01001101",
        223 => "01001100",
        222 => "01001011",
        221 => "01001010",
        220 => "01001001",
        219 => "01001000",
        218 => "01000111",
        217 => "01000111",
        216 => "01000110",
        215 => "01000101",
        214 => "01000101",
        213 => "01000100",
        212 => "01000011",
        211 => "01000011",
        210 => "01000010",
        209 => "01000001",
        208 => "01000001",
        207 => "01000000",
        206 => "01000000",
        205 => "00111111",
        204 => "00111110",
        203 => "00111110",
        202 => "00111101",
        201 => "00111101",
        200 => "00111100",
        199 => "00111100",
        198 => "00111011",
        197 => "00111011",
        196 => "00111010",
        195 => "00111010",
        194 => "00111010",
        193 => "00111001",
        192 => "00111001",
        191 => "00111000",
        190 => "00111000",
        189 => "00110111",
        188 => "00110111",
        187 => "00110110",
        186 => "00110110",
        185 => "00110110",
        184 => "00110101",
        183 => "00110101",
        182 => "00110100",
        181 => "00110100",
        180 => "00110100",
        179 => "00110011",
        178 => "00110011",
        177 => "00110010",
        176 => "00110010",
        175 => "00110010",
        174 => "00110001",
        173 => "00110001",
        172 => "00110000",
        171 => "00110000",
        170 => "00110000",
        169 => "00101111",
        168 => "00101111",
        167 => "00101111",
        166 => "00101110",
        165 => "00101110",
        164 => "00101101",
        163 => "00101101",
        162 => "00101101",
        161 => "00101100",
        160 => "00101100",
        159 => "00101100",
        158 => "00101011",
        157 => "00101011",
        156 => "00101011",
        155 => "00101010",
        154 => "00101010",
        153 => "00101010",
        152 => "00101001",
        151 => "00101001",
        150 => "00101001",
        149 => "00101000",
        148 => "00101000",
        147 => "00101000",
        146 => "00100111",
        145 => "00100111",
        144 => "00100111",
        143 => "00100110",
        142 => "00100110",
        141 => "00100110",
        140 => "00100101",
        139 => "00100101",
        138 => "00100101",
        137 => "00100101",
        136 => "00100100",
        135 => "00100100",
        134 => "00100100",
        133 => "00100011",
        132 => "00100011",
        131 => "00100011",
        130 => "00100010",
        129 => "00100010",
        128 => "00100010",
        127 => "00100010",
        126 => "00100001",
        125 => "00100001",
        124 => "00100001",
        123 => "00100000",
        122 => "00100000",
        121 => "00100000",
        120 => "00011111",
        119 => "00011111",
        118 => "00011111",
        117 => "00011111",
        116 => "00011110",
        115 => "00011110",
        114 => "00011110",
        113 => "00011101",
        112 => "00011101",
        111 => "00011101",
        110 => "00011101",
        109 => "00011100",
        108 => "00011100",
        107 => "00011100",
        106 => "00011011",
        105 => "00011011",
        104 => "00011011",
        103 => "00011011",
        102 => "00011010",
        101 => "00011010",
        100 => "00011010",
        99 => "00011001",
        98 => "00011001",
        97 => "00011001",
        96 => "00011001",
        95 => "00011000",
        94 => "00011000",
        93 => "00011000",
        92 => "00011000",
        91 => "00010111",
        90 => "00010111",
        89 => "00010111",
        88 => "00010110",
        87 => "00010110",
        86 => "00010110",
        85 => "00010110",
        84 => "00010101",
        83 => "00010101",
        82 => "00010101",
        81 => "00010101",
        80 => "00010100",
        79 => "00010100",
        78 => "00010100",
        77 => "00010100",
        76 => "00010011",
        75 => "00010011",
        74 => "00010011",
        73 => "00010011",
        72 => "00010010",
        71 => "00010010",
        70 => "00010010",
        69 => "00010001",
        68 => "00010001",
        67 => "00010001",
        66 => "00010001",
        65 => "00010000",
        64 => "00010000",
        63 => "00010000",
        62 => "00010000",
        61 => "00001111",
        60 => "00001111",
        59 => "00001111",
        58 => "00001111",
        57 => "00001110",
        56 => "00001110",
        55 => "00001110",
        54 => "00001110",
        53 => "00001101",
        52 => "00001101",
        51 => "00001101",
        50 => "00001101",
        49 => "00001100",
        48 => "00001100",
        47 => "00001100",
        46 => "00001100",
        45 => "00001011",
        44 => "00001011",
        43 => "00001011",
        42 => "00001011",
        41 => "00001010",
        40 => "00001010",
        39 => "00001010",
        38 => "00001010",
        37 => "00001001",
        36 => "00001001",
        35 => "00001001",
        34 => "00001001",
        33 => "00001000",
        32 => "00001000",
        31 => "00001000",
        30 => "00000111",
        29 => "00000111",
        28 => "00000111",
        27 => "00000111",
        26 => "00000110",
        25 => "00000110",
        24 => "00000110",
        23 => "00000110",
        22 => "00000101",
        21 => "00000101",
        20 => "00000101",
        19 => "00000101",
        18 => "00000100",
        17 => "00000100",
        16 => "00000100",
        15 => "00000100",
        14 => "00000011",
        13 => "00000011",
        12 => "00000011",
        11 => "00000011",
        10 => "00000010",
        9 => "00000010",
        8 => "00000010",
        7 => "00000010",
        6 => "00000001",
        5 => "00000001",
        4 => "00000001",
        3 => "00000001",
        2 => "00000000",
        1 => "00000000",
        0 => "00000000"
    );



begin
    process(raw_in)
    begin
        if signal_bit = '0' then  -- Substitua ":" por "then" e use "=" ao invés de "=="
            -- Converte a entrada para inteiro e seleciona o valor da tabela
            angle_out <= angle_table(to_integer(unsigned(raw_in)));
        else
            angle_out <= negative_angle_table(to_integer(unsigned(raw_in)));
            --angle_out <= "01010101";
        end if;  -- Encerramento do bloco if
    end process;
end architecture rtl;

