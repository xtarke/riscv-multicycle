library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.M_types.all;

entity M is
	port(
		CLOCK :in std_logic;
		M_data : in M_data_t;		
		dataOut  : out std_logic_vector(31 downto 0)
	);
end entity;

architecture RTL of M is
	-------------------------------------------------------------------	


	signal mul_logic_vector: Signed(63 downto 0);
	signal mulu_logic_vector: Unsigned(63 downto 0);
	
	signal div_logic_vector: Signed(31 downto 0);
	signal divu_logic_vector: Unsigned(31 downto 0);
	
	signal rem_logic_vector: Signed(31 downto 0);
	signal remu_logic_vector: Unsigned(31 downto 0);

begin
	--===============================================================--

	mul_logic_vector <= M_data.a*M_data.b;
	mulu_logic_vector <= Unsigned(M_data.a)*Unsigned(M_data.b);

	div_logic_vector <= M_data.a/M_data.b;
	divu_logic_vector <= Unsigned(M_data.a)/Unsigned(M_data.b);
	
	rem_logic_vector <= M_data.a mod M_data.b;  
	remu_logic_vector <= Unsigned(M_data.a) mod Unsigned(M_data.b);

	ula_op : with M_data.code select
		dataOut <=	Std_logic_vector(mul_logic_vector(31 downto 0)) when M_MUL,
					Std_logic_vector(mul_logic_vector(63 downto 32)) when M_MULH,

					Std_logic_vector(mulu_logic_vector(63 downto 32)) when M_MULHU,
					Std_logic_vector(mulu_logic_vector(63 downto 32)) when M_MULHSU,

					Std_logic_vector(div_logic_vector) when M_DIV,
					Std_logic_vector(divu_logic_vector) when M_DIVU,
					
					Std_logic_vector(rem_logic_vector) when M_REM,
					Std_logic_vector(remu_logic_vector) when M_REMU,
			        (others => '0') when others;

end architecture;