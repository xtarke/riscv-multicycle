-------------------------------------------------------------------
-- Name        : de0_lite.vhd
-- Author      : 
-- Version     : 0.1
-- Copyright   : Departamento de Eletrônica, Florianópolis, IFSC
-- Description : Projeto base DE10-Lite
-------------------------------------------------------------------
LIBRARY ieee;
USE IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;
-- Utilização das funções de my_package
use work.logica7.all;

entity de10_lite is 
	port (
		---------- CLOCK ----------
		ADC_CLK_10:	in std_logic;
		MAX10_CLK1_50: in std_logic;
		MAX10_CLK2_50: in std_logic;
		
		----------- SDRAM ------------
		DRAM_ADDR: out std_logic_vector (12 downto 0);
		DRAM_BA: out std_logic_vector (1 downto 0);
		DRAM_CAS_N: out std_logic;
		DRAM_CKE: out std_logic;
		DRAM_CLK: out std_logic;
		DRAM_CS_N: out std_logic;		
		DRAM_DQ: inout std_logic_vector(15 downto 0);
		DRAM_LDQM: out std_logic;
		DRAM_RAS_N: out std_logic;
		DRAM_UDQM: out std_logic;
		DRAM_WE_N: out std_logic;
		
		----------- SEG7 ------------
		HEX0: out std_logic_vector(7 downto 0);
		HEX1: out std_logic_vector(7 downto 0);
		HEX2: out std_logic_vector(7 downto 0);
		HEX3: out std_logic_vector(7 downto 0);
		HEX4: out std_logic_vector(7 downto 0);
		HEX5: out std_logic_vector(7 downto 0);

		----------- KEY ------------
		KEY: in std_logic_vector(1 downto 0);

		----------- LED ------------
		LEDR: out std_logic_vector(9 downto 0);

		----------- SW ------------
		SW: in std_logic_vector(9 downto 0);

		----------- VGA ------------
		VGA_B: out std_logic_vector(3 downto 0);
		VGA_G: out std_logic_vector(3 downto 0);
		VGA_HS: out std_logic;
		VGA_R: out std_logic_vector(3 downto 0);
		VGA_VS: out std_logic;
	
		----------- Accelerometer ------------
		GSENSOR_CS_N: out std_logic;
		GSENSOR_INT: in std_logic_vector(2 downto 1);
		GSENSOR_SCLK: out std_logic;
		GSENSOR_SDI: inout std_logic;
		GSENSOR_SDO: inout std_logic;
	
		----------- Arduino ------------
		ARDUINO_IO: inout std_logic_vector(15 downto 0);
		ARDUINO_RESET_N: inout std_logic
	);
end entity;


architecture rtl of de10_lite is


	signal frequencia: unsigned(31 downto 0);


begin
	

	   
	   encoder:entity work.encoder
	       port map(
	           clk           => MAX10_CLK1_50,
	           aclr_n        => SW(0),
	           select_time   => SW(4 downto 2),
	           encoder_pulse => SW(1),
	           frequency     => frequencia
	       );
	   
	       display0:entity work.seven_segment_cntrl
            port map(
                input => frequencia(3 downto 0),
                segs  => HEX0
            );
            
            display1:entity work.seven_segment_cntrl
            port map(
                input => frequencia(7 downto 4),
                segs  => HEX1
            );
	    
           display2:entity work.seven_segment_cntrl
            port map(
                input => frequencia(11 downto 8),
                segs  => HEX2
            );
           display3:entity work.seven_segment_cntrl
            port map(
                input => frequencia(15 downto 12),
                segs  => HEX3
            );
            
            display4:entity work.seven_segment_cntrl
            port map(
                input => frequencia(19 downto 16),
                segs  => HEX4
            );
           display5:entity work.seven_segment_cntrl
            port map(
                input => frequencia(23 downto 20),
                segs  => HEX5
            );
end;

