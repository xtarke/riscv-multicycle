
module rotacao (
	source);	

	output	[31:0]	source;
endmodule
