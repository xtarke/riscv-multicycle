library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity filename is
    port(
        clk : in std_logic;
        rst : in std_logic
    );
end entity filename;

architecture RTL of filename is
    
begin

end architecture RTL;
