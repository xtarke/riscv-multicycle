
module probes (
	source,
	probe);	

	output	[19:0]	source;
	input	[19:0]	probe;
endmodule
