-------------------------------------------------------
--! @file    heaviside.vhd
--! @author  Leonardo Benitez
--! @date    2021-11-02
--! @version 0.1
--! @brief   Decoder for seven segments display; 
--!          Leds are active in 0
-------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity heaviside is
    port (
        input:       in  std_logic_vector(7 downto 0);
        output:        out std_logic_vector(7 downto 0)
    );
end entity heaviside;

architecture rtl of heaviside is
begin
	process (input)
	begin
		case input is				
		when "10000000" => output <= "00000000";  -- -128
		when "10000001" => output <= "00000000";  -- -127
		when "10000010" => output <= "00000000";  -- -126
		when "10000011" => output <= "00000000";  -- -125
		when "10000100" => output <= "00000000";  -- -124
		when "10000101" => output <= "00000000";  -- -123
		when "10000110" => output <= "00000000";  -- -122
		when "10000111" => output <= "00000000";  -- -121
		when "10001000" => output <= "00000000";  -- -120
		when "10001001" => output <= "00000000";  -- -119
		when "10001010" => output <= "00000000";  -- -118
		when "10001011" => output <= "00000000";  -- -117
		when "10001100" => output <= "00000000";  -- -116
		when "10001101" => output <= "00000000";  -- -115
		when "10001110" => output <= "00000000";  -- -114
		when "10001111" => output <= "00000000";  -- -113
		when "10010000" => output <= "00000000";  -- -112
		when "10010001" => output <= "00000000";  -- -111
		when "10010010" => output <= "00000000";  -- -110
		when "10010011" => output <= "00000000";  -- -109
		when "10010100" => output <= "00000000";  -- -108
		when "10010101" => output <= "00000000";  -- -107
		when "10010110" => output <= "00000000";  -- -106
		when "10010111" => output <= "00000000";  -- -105
		when "10011000" => output <= "00000000";  -- -104
		when "10011001" => output <= "00000000";  -- -103
		when "10011010" => output <= "00000000";  -- -102
		when "10011011" => output <= "00000000";  -- -101
		when "10011100" => output <= "00000000";  -- -100
		when "10011101" => output <= "00000000";  -- -99
		when "10011110" => output <= "00000000";  -- -98
		when "10011111" => output <= "00000000";  -- -97
		when "10100000" => output <= "00000000";  -- -96
		when "10100001" => output <= "00000000";  -- -95
		when "10100010" => output <= "00000000";  -- -94
		when "10100011" => output <= "00000000";  -- -93
		when "10100100" => output <= "00000000";  -- -92
		when "10100101" => output <= "00000000";  -- -91
		when "10100110" => output <= "00000000";  -- -90
		when "10100111" => output <= "00000000";  -- -89
		when "10101000" => output <= "00000000";  -- -88
		when "10101001" => output <= "00000000";  -- -87
		when "10101010" => output <= "00000000";  -- -86
		when "10101011" => output <= "00000000";  -- -85
		when "10101100" => output <= "00000000";  -- -84
		when "10101101" => output <= "00000000";  -- -83
		when "10101110" => output <= "00000000";  -- -82
		when "10101111" => output <= "00000000";  -- -81
		when "10110000" => output <= "00000000";  -- -80
		when "10110001" => output <= "00000000";  -- -79
		when "10110010" => output <= "00000000";  -- -78
		when "10110011" => output <= "00000000";  -- -77
		when "10110100" => output <= "00000000";  -- -76
		when "10110101" => output <= "00000000";  -- -75
		when "10110110" => output <= "00000000";  -- -74
		when "10110111" => output <= "00000000";  -- -73
		when "10111000" => output <= "00000000";  -- -72
		when "10111001" => output <= "00000000";  -- -71
		when "10111010" => output <= "00000000";  -- -70
		when "10111011" => output <= "00000000";  -- -69
		when "10111100" => output <= "00000000";  -- -68
		when "10111101" => output <= "00000000";  -- -67
		when "10111110" => output <= "00000000";  -- -66
		when "10111111" => output <= "00000000";  -- -65
		when "11000000" => output <= "00000000";  -- -64
		when "11000001" => output <= "00000000";  -- -63
		when "11000010" => output <= "00000000";  -- -62
		when "11000011" => output <= "00000000";  -- -61
		when "11000100" => output <= "00000000";  -- -60
		when "11000101" => output <= "00000000";  -- -59
		when "11000110" => output <= "00000000";  -- -58
		when "11000111" => output <= "00000000";  -- -57
		when "11001000" => output <= "00000000";  -- -56
		when "11001001" => output <= "00000000";  -- -55
		when "11001010" => output <= "00000000";  -- -54
		when "11001011" => output <= "00000000";  -- -53
		when "11001100" => output <= "00000000";  -- -52
		when "11001101" => output <= "00000000";  -- -51
		when "11001110" => output <= "00000000";  -- -50
		when "11001111" => output <= "00000000";  -- -49
		when "11010000" => output <= "00000000";  -- -48
		when "11010001" => output <= "00000000";  -- -47
		when "11010010" => output <= "00000000";  -- -46
		when "11010011" => output <= "00000000";  -- -45
		when "11010100" => output <= "00000000";  -- -44
		when "11010101" => output <= "00000000";  -- -43
		when "11010110" => output <= "00000000";  -- -42
		when "11010111" => output <= "00000000";  -- -41
		when "11011000" => output <= "00000000";  -- -40
		when "11011001" => output <= "00000000";  -- -39
		when "11011010" => output <= "00000000";  -- -38
		when "11011011" => output <= "00000000";  -- -37
		when "11011100" => output <= "00000000";  -- -36
		when "11011101" => output <= "00000000";  -- -35
		when "11011110" => output <= "00000000";  -- -34
		when "11011111" => output <= "00000000";  -- -33
		when "11100000" => output <= "00000000";  -- -32
		when "11100001" => output <= "00000000";  -- -31
		when "11100010" => output <= "00000000";  -- -30
		when "11100011" => output <= "00000000";  -- -29
		when "11100100" => output <= "00000000";  -- -28
		when "11100101" => output <= "00000000";  -- -27
		when "11100110" => output <= "00000000";  -- -26
		when "11100111" => output <= "00000000";  -- -25
		when "11101000" => output <= "00000000";  -- -24
		when "11101001" => output <= "00000000";  -- -23
		when "11101010" => output <= "00000000";  -- -22
		when "11101011" => output <= "00000000";  -- -21
		when "11101100" => output <= "00000000";  -- -20
		when "11101101" => output <= "00000000";  -- -19
		when "11101110" => output <= "00000000";  -- -18
		when "11101111" => output <= "00000000";  -- -17
		when "11110000" => output <= "00000000";  -- -16
		when "11110001" => output <= "00000000";  -- -15
		when "11110010" => output <= "00000000";  -- -14
		when "11110011" => output <= "00000000";  -- -13
		when "11110100" => output <= "00000000";  -- -12
		when "11110101" => output <= "00000000";  -- -11
		when "11110110" => output <= "00000000";  -- -10
		when "11110111" => output <= "00000000";  -- -9
		when "11111000" => output <= "00000000";  -- -8
		when "11111001" => output <= "00000000";  -- -7
		when "11111010" => output <= "00000000";  -- -6
		when "11111011" => output <= "00000000";  -- -5
		when "11111100" => output <= "00000000";  -- -4
		when "11111101" => output <= "00000000";  -- -3
		when "11111110" => output <= "00000000";  -- -2
		when "11111111" => output <= "00000000";  -- -1
		when "00000000" => output <= "00000000";  -- 0
		when "00000001" => output <= "01111111";  -- 1
		when "00000010" => output <= "01111111";  -- 2
		when "00000011" => output <= "01111111";  -- 3
		when "00000100" => output <= "01111111";  -- 4
		when "00000101" => output <= "01111111";  -- 5
		when "00000110" => output <= "01111111";  -- 6
		when "00000111" => output <= "01111111";  -- 7
		when "00001000" => output <= "01111111";  -- 8
		when "00001001" => output <= "01111111";  -- 9
		when "00001010" => output <= "01111111";  -- 10
		when "00001011" => output <= "01111111";  -- 11
		when "00001100" => output <= "01111111";  -- 12
		when "00001101" => output <= "01111111";  -- 13
		when "00001110" => output <= "01111111";  -- 14
		when "00001111" => output <= "01111111";  -- 15
		when "00010000" => output <= "01111111";  -- 16
		when "00010001" => output <= "01111111";  -- 17
		when "00010010" => output <= "01111111";  -- 18
		when "00010011" => output <= "01111111";  -- 19
		when "00010100" => output <= "01111111";  -- 20
		when "00010101" => output <= "01111111";  -- 21
		when "00010110" => output <= "01111111";  -- 22
		when "00010111" => output <= "01111111";  -- 23
		when "00011000" => output <= "01111111";  -- 24
		when "00011001" => output <= "01111111";  -- 25
		when "00011010" => output <= "01111111";  -- 26
		when "00011011" => output <= "01111111";  -- 27
		when "00011100" => output <= "01111111";  -- 28
		when "00011101" => output <= "01111111";  -- 29
		when "00011110" => output <= "01111111";  -- 30
		when "00011111" => output <= "01111111";  -- 31
		when "00100000" => output <= "01111111";  -- 32
		when "00100001" => output <= "01111111";  -- 33
		when "00100010" => output <= "01111111";  -- 34
		when "00100011" => output <= "01111111";  -- 35
		when "00100100" => output <= "01111111";  -- 36
		when "00100101" => output <= "01111111";  -- 37
		when "00100110" => output <= "01111111";  -- 38
		when "00100111" => output <= "01111111";  -- 39
		when "00101000" => output <= "01111111";  -- 40
		when "00101001" => output <= "01111111";  -- 41
		when "00101010" => output <= "01111111";  -- 42
		when "00101011" => output <= "01111111";  -- 43
		when "00101100" => output <= "01111111";  -- 44
		when "00101101" => output <= "01111111";  -- 45
		when "00101110" => output <= "01111111";  -- 46
		when "00101111" => output <= "01111111";  -- 47
		when "00110000" => output <= "01111111";  -- 48
		when "00110001" => output <= "01111111";  -- 49
		when "00110010" => output <= "01111111";  -- 50
		when "00110011" => output <= "01111111";  -- 51
		when "00110100" => output <= "01111111";  -- 52
		when "00110101" => output <= "01111111";  -- 53
		when "00110110" => output <= "01111111";  -- 54
		when "00110111" => output <= "01111111";  -- 55
		when "00111000" => output <= "01111111";  -- 56
		when "00111001" => output <= "01111111";  -- 57
		when "00111010" => output <= "01111111";  -- 58
		when "00111011" => output <= "01111111";  -- 59
		when "00111100" => output <= "01111111";  -- 60
		when "00111101" => output <= "01111111";  -- 61
		when "00111110" => output <= "01111111";  -- 62
		when "00111111" => output <= "01111111";  -- 63
		when "01000000" => output <= "01111111";  -- 64
		when "01000001" => output <= "01111111";  -- 65
		when "01000010" => output <= "01111111";  -- 66
		when "01000011" => output <= "01111111";  -- 67
		when "01000100" => output <= "01111111";  -- 68
		when "01000101" => output <= "01111111";  -- 69
		when "01000110" => output <= "01111111";  -- 70
		when "01000111" => output <= "01111111";  -- 71
		when "01001000" => output <= "01111111";  -- 72
		when "01001001" => output <= "01111111";  -- 73
		when "01001010" => output <= "01111111";  -- 74
		when "01001011" => output <= "01111111";  -- 75
		when "01001100" => output <= "01111111";  -- 76
		when "01001101" => output <= "01111111";  -- 77
		when "01001110" => output <= "01111111";  -- 78
		when "01001111" => output <= "01111111";  -- 79
		when "01010000" => output <= "01111111";  -- 80
		when "01010001" => output <= "01111111";  -- 81
		when "01010010" => output <= "01111111";  -- 82
		when "01010011" => output <= "01111111";  -- 83
		when "01010100" => output <= "01111111";  -- 84
		when "01010101" => output <= "01111111";  -- 85
		when "01010110" => output <= "01111111";  -- 86
		when "01010111" => output <= "01111111";  -- 87
		when "01011000" => output <= "01111111";  -- 88
		when "01011001" => output <= "01111111";  -- 89
		when "01011010" => output <= "01111111";  -- 90
		when "01011011" => output <= "01111111";  -- 91
		when "01011100" => output <= "01111111";  -- 92
		when "01011101" => output <= "01111111";  -- 93
		when "01011110" => output <= "01111111";  -- 94
		when "01011111" => output <= "01111111";  -- 95
		when "01100000" => output <= "01111111";  -- 96
		when "01100001" => output <= "01111111";  -- 97
		when "01100010" => output <= "01111111";  -- 98
		when "01100011" => output <= "01111111";  -- 99
		when "01100100" => output <= "01111111";  -- 100
		when "01100101" => output <= "01111111";  -- 101
		when "01100110" => output <= "01111111";  -- 102
		when "01100111" => output <= "01111111";  -- 103
		when "01101000" => output <= "01111111";  -- 104
		when "01101001" => output <= "01111111";  -- 105
		when "01101010" => output <= "01111111";  -- 106
		when "01101011" => output <= "01111111";  -- 107
		when "01101100" => output <= "01111111";  -- 108
		when "01101101" => output <= "01111111";  -- 109
		when "01101110" => output <= "01111111";  -- 110
		when "01101111" => output <= "01111111";  -- 111
		when "01110000" => output <= "01111111";  -- 112
		when "01110001" => output <= "01111111";  -- 113
		when "01110010" => output <= "01111111";  -- 114
		when "01110011" => output <= "01111111";  -- 115
		when "01110100" => output <= "01111111";  -- 116
		when "01110101" => output <= "01111111";  -- 117
		when "01110110" => output <= "01111111";  -- 118
		when "01110111" => output <= "01111111";  -- 119
		when "01111000" => output <= "01111111";  -- 120
		when "01111001" => output <= "01111111";  -- 121
		when "01111010" => output <= "01111111";  -- 122
		when "01111011" => output <= "01111111";  -- 123
		when "01111100" => output <= "01111111";  -- 124
		when "01111101" => output <= "01111111";  -- 125
		when "01111110" => output <= "01111111";  -- 126
		when others => output <= "01111111";  -- 127
		end case;
	end process;
end architecture rtl;